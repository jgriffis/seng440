----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:23:08 08/18/2013 
-- Design Name: 
-- Module Name:    lookup - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity lookup is
	Port (
		argument : in STD_LOGIC_VECTOR (6 downto 0);
		symbol : out STD_LOGIC_VECTOR (3 downto 0);
		code_length : out STD_LOGIC_VECTOR (3 downto 0)
	);
end lookup;

architecture Behavioral of lookup is

	type lut is array (0 to 127) of STD_LOGIC_VECTOR(7 downto 0);
	constant hd_lut  : lut  := 
	( 0 => "10110011",
	  1 => "10110011",
	  2 => "10110011",
	  3 => "10110011",
	  4 => "10110011",
	  5 => "10110011",
	  6 => "10110011",
	  7 => "10110011",
	  8 => "10110011",
	  9 => "10110011",
	 10 => "10110011",
	 11 => "10110011",
	 12 => "10110011",
	 13 => "10110011",
	 14 => "10110011",
	 15 => "10110011",
	 16 => "11000011",
	 17 => "11000011",
	 18 => "11000011",
	 19 => "11000011",
	 20 => "11000011",
	 21 => "11000011",
	 22 => "11000011",
	 23 => "11000011",
	 24 => "11000011",
	 25 => "11000011",
	 26 => "11000011",
	 27 => "11000011",
	 28 => "11000011",
	 29 => "11000011",
	 30 => "11000011",
	 31 => "11000011",
	 32 => "01110100",
	 33 => "01110100",
	 34 => "01110100",
	 35 => "01110100",
	 36 => "01110100",
	 37 => "01110100",
	 38 => "01110100",
	 39 => "01110100",
	 40 => "01100101",
	 41 => "01100101",
	 42 => "01100101",
	 43 => "01100101",
	 44 => "01010101",
	 45 => "01010101",
	 46 => "01010101",
	 47 => "01010101",
	 48 => "10000100",
	 49 => "10000100",
	 50 => "10000100",
	 51 => "10000100",
	 52 => "10000100",
	 53 => "10000100",
	 54 => "10000100",
	 55 => "10000100",
	 56 => "10010100",
	 57 => "10010100",
	 58 => "10010100",
	 59 => "10010100",
	 60 => "10010100",
	 61 => "10010100",
	 62 => "10010100",
	 63 => "10010100",
	 64 => "11010011",
	 65 => "11010011",
	 66 => "11010011",
	 67 => "11010011",
	 68 => "11010011",
	 69 => "11010011",
	 70 => "11010011",
	 71 => "11010011",
	 72 => "11010011",
	 73 => "11010011",
	 74 => "11010011",
	 75 => "11010011",
	 76 => "11010011",
	 77 => "11010011",
	 78 => "11010011",
	 79 => "11010011",
	 80 => "11100011",
	 81 => "11100011",
	 82 => "11100011",
	 83 => "11100011",
	 84 => "11100011",
	 85 => "11100011",
	 86 => "11100011",
	 87 => "11100011",
	 88 => "11100011",
	 89 => "11100011",
	 90 => "11100011",
	 91 => "11100011",
	 92 => "11100011",
	 93 => "11100011",
	 94 => "11100011",
	 95 => "11100011",
	 96 => "10100100",
	 97 => "10100100",
	 98 => "10100100",
	 99 => "10100100",
	100 => "10100100",
	101 => "10100100",
	102 => "10100100",
	103 => "10100100",
	104 => "01000110",
	105 => "01000110",
	106 => "00110110",
	107 => "00110110",
	108 => "00000111",
	109 => "00010111",
	110 => "00100110",
	111 => "00100110",
	112 => "11110011",
	113 => "11110011",
	114 => "11110011",
	115 => "11110011",
	116 => "11110011",
	117 => "11110011",
	118 => "11110011",
	119 => "11110011",
	120 => "11110011",
	121 => "11110011",
	122 => "11110011",
	123 => "11110011",
	124 => "11110011",
	125 => "11110011",
	126 => "11110011",
	127 => "11110011");

begin

	process (argument)
	begin
		symbol 		<= hd_lut(to_integer(unsigned(argument))) (7 downto 4);
		code_length <= hd_lut(to_integer(unsigned(argument))) (3 downto 0);
	end process;

end Behavioral;

